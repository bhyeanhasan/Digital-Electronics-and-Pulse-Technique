* C:\Users\NoYoN\Desktop\Digital-Electronics-and-Pulse-Technique\mid.sch

* Schematics Version 9.1 - Web Update 1
* Thu Aug 03 16:46:25 2023



** Analysis setup **
.tran 0ns 100m
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "mid.net"
.INC "mid.als"


.probe


.END
